* This file contains all the subcircuits to be used in SRAM256.cir

***** long channel VTP = -0.9, VTN = 0.8 *****
*.include modelcard/1um.pm
*.param supply = 5
*.param ll = 1u

****** 50nm models***


.include 50nm.pm
.param supply =1

.param lambda=25nm
.param ll='2*lambda'

****** 16nm low power models***
*.include ./modelcard/PTM_LP/16nm.pm
*.param supply =0.9
*.param ll=16nm

****** 16nm high peformance models***
*.include ./modelcard/PTM_HP/16nm.pm
*.param supply =0.7
*.param ll=16nm


.subckt wire iot iof len=10 wid=10
.param rr=0.4
.param cc = '100e-15'
rt iot iof 'rr*len*50/(wid)'
cf iof  0  'cc*len*wid*50/1e6'

.ends

.subckt wire_dual lt rt lf rf len=10 wid=10
Xt lt rt wire len='len' wid='wid'
Xf lf rf wire len='len' wid='wid'
.ends

.subckt nn d g s  ww=100
mnfet d g s 0 nmos L=ll w='ww*ll'
.ends

.subckt pp d g s   ww=100
mpfet d g s vdd pmos L=ll w='ww*ll'
.ends


.subckt inv out inn size=30 beta=2
XPP out inn vdd pp ww='size*beta/(beta+1)'
XNN out inn gnd nn ww='size/(beta+1)'
.ends

.subckt nnd2 out in1 in0 size=30 beta=2
Xap0 out in0 vdd pp ww='beta*size/(beta+2)'
Xap1 out in1 vdd pp ww='beta*size/(beta+2)'
Xan0 out in0 nng nn ww='2*size/(beta+2)'
Xan1 nng in1 0   nn ww='2*size/(beta+2)'
.ends nnd2

.subckt nor2 out in1 in0 size=30 beta=2
Xap0 ppi in0 vdd pp ww='2*beta*size/(2*beta+1)'
Xap1 out in1 ppi pp ww='2*beta*size/(2*beta+1)'
Xan0 out in0 0 nn ww='1*size/(2*beta+1)'
Xan1 out in1 0   nn ww='1*size/(2*beta+1)'
.ends nor2

.subckt latch out inn clk clb size=15 beta=2
Xn inn clk qin nn ww='5'
Xp inn clb qin pp ww='10'

Xfp qin ggg vdd pp ww='5'
Xfn qin ggg gnd nn ww='5'

Xi ggg qin     inv size='size'
Xo out ggg     inv size='3*size'
.ends latch

.subckt flop qqq ddd clk
Xinve clb clk inv
Xflip int ddd clb clk latch
Xflop qqq int clk clb latch
.ends flop

.subckt reg8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 clk
x7 ot7 in7 clk flop
x6 ot6 in6 clk flop
x5 ot5 in5 clk flop
x4 ot4 in4 clk flop
x3 ot3 in3 clk flop
x2 ot2 in2 clk flop
x1 ot1 in1 clk flop
x0 ot0 in0 clk flop
.ends reg8

.subckt dat1 out period=1ns start=1ns sz=50 total=5 duty=3
V0 j0  0  PULSE('supply' 0 'start' 10p 10p 'duty*period-10ps' 'total*period')
x7 out j0 inv size='sz'
.ends dat1

*generates different data stream on all eight channels, buffered output
.subckt dat8 o7 o6 o5 o4 o3 o2 o1 o0 per=1ns start=1ns size=50
V0 j0  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' 'per')
V1 j1  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '2*per')
V2 j2  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '3*per')
V3 j3  0  PULSE(0 'supply' 'start' 10p 10p '0.5*per-10ps' '4*per')
V4 j4  0  PULSE('supply' 0 'start' 10p 10p '0.5*per-10ps' '1*per')
V5 j5  0  PULSE('supply' 0 'start' 10p 10p '1*per-10ps' '2*per')
V6 j6  0  PULSE('supply' 0 'start' 10p 10p '1.5*per-10ps' '3*per')
V7 j7  0  PULSE('supply' 0 'start' 10p 10p '2*per-10ps' '4*per')
xb o7 o6 o5 o4 o3 o2 o1 o0 j7 j6 j5 j4 j3 j2 j1 j0 buf8 sz='size'
.ends dat8

.subckt buf8 ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0 in7 in6 in5 in4 in3 in2 in1 in0 sz=100
x7 ot7 in7 inv size='sz'
x6 ot6 in6 inv size='sz'
x5 ot5 in5 inv size='sz'
x4 ot4 in4 inv size='sz'
x3 ot3 in3 inv size='sz'
x2 ot2 in2 inv size='sz'
x1 ot1 in1 inv size='sz'
x0 ot0 in0 inv size='sz'
.ends buf8


.subckt nnd3 out in2 in1 in0 size=20 beta=2
Xp0 out in0 vdd pp ww='beta*size/(beta+3)'
Xp1 out in1 vdd pp ww='beta*size/(beta+3)'
Xp2 out in2 vdd pp ww='beta*size/(beta+3)'
Xn0 out in0 nn0 nn ww='3*size/(beta+3)'
Xn1 nn0 in1 nn1 nn ww='3*size/(beta+3)'
Xn2 nn1 in2 gnd nn ww='3*size/(beta+3)'
.ends

.subckt senseAmp ot1 ot0 in1 in0 eva size=40
Xn0 ot0 in0 ot1 eva nnd3 size ='size'
Xn1 ot1 in1 ot0 eva nnd3 size ='size'
.ends senseAmp

*can improve this at the Xnd5 area
.subckt decModel cho din clk sz=100
Xi1  nn1 din     inv  size='sz'
Xnd2 nn2 nn1 vdd nnd2 size='2*sz'
xdu2 dd1 nn1 gnd nnd2 size='2*sz'
xnr3 nn3 nn2 gnd nor2 size='5*sz'
xdu3 dd2 nn2 vdd nor2 size='5*sz*3'
Xnd4 nn4 nn3 vdd nnd2 size='2*sz'
xdu4 dd3 nn3 gnd nnd2 size='30sz*1'
Xnd5 nn5 nn4 clk nnd2 size='2*sz'
Xin6 cho nn5     inv  size='sz'
.ends



.subckt write_buffer btt bff dii rwt clk adr
Xi1   nn1 clk          inv
Xi2   nn2 nn1          inv
Xi3   trg nn2          inv
Xnr1  nn3 trg rwt adr  nor3
Xnn1  nn4 nn3 gnd      nn
Xnn2  btt dii nn4      nn
Xpp1  btt nn3 vdd      pp
Xi4   nn5 dii          inv
Xnn3  nn6 nn3 gnd      nn
Xnn4  bff nn5 nn6      nn
Xpp2  bff nn3 vdd      pp
.ends write_buffer



.subckt write1 btt bff dii rwt clk sz=10
Xi1   nn1 clk     inv
Xi2   nn2 nn1     inv size='50'
Xi3   trg nn2     inv
Xnr1  nn3 trg rwt nor2 size='sz*2'
Xpp1  btt nn3 vdd pp   size='sz'
Xnn1  btt nn3 nn4 nn   size='sz*3'
Xnn2  nn4 dii gnd nn   size='sz*3'
Xi4   nn5 dii     inv  size='sz'
Xpp2  bff nn3 vdd pp   size='sz'
xnn3  bff nn3 nn6 nn   size='sz*3'
Xnn4  nn6 nn5 gnd nn   size='sz*3'
.ends write1



.subckt read1 btt bff dot rwt clk
Xnd1  nn1 rwt clk         nnd2     size='10'
Xi1   trg nn1             inv      size='20'
Xsns1 tru fal btt bff trg senseAmp size='50'
Xi2   nn2 tru             inv      size='20'
Xi3   nn3 fal             inv      size='20'
Xi4   nn4 nn3             inv      size='20'
Xpp1  dot nn4 vdd         pp	   ww='20'
Xnn1  dot nn2 gnd         nn       ww='10'
Xi5   dot nn5             inv      size='10'
Xi6   nn5 dot             inv
.ends read1


.subckt readSub btt bff set rst sel rdw clk
Xsns1 set rst btt bff trg senseAmp sz='50'
Xnnd3 trgn sel clk rdw    nnd3
X0    trg trgn            inv size='150'

.ends readSub


.subckt readcollect dot st3 rs3 st2 rs2 st1 rs1 st0 rs0
Xset0 aa0 st3 st2 nnd2
Xset1 aa1 st1 st0 nnd2
X0    hi0 aa0     inv
X1    hi1 aa1     inv
Xrs0  lo1 rs3 rs2 nnd2
Xrs1  lo0 rs1 rs0 nnd2
Xp0   dot hi0 vdd pp
Xp1   dot hi1 vdd pp
Xn0   dot lo1 gnd nn
Xn1   dot lo0 gnd nn
X2    nnn dot     inv size='5' beta=1
X3    dot nnn     inv size='5' beta=1
.ends readcollect


.subckt subblock set rst add din rdw clk lw=2368 wirew=10
Xwr bt1 bf1 din rdw clk         writeSub
Xw1 bt1 btt bf1 bff             wire_dual len'lw' wid'wirew'
Xmd btt bff                     memLoad number=31
Xla btt bff clk                 mem1
Xrd btt bff set rst bdd rdw clk readSub
.ends subblock

.subckt mem1 bff btt wl
Xn1  Qn  Q  gnd nn ww='5'
Xp2  Qn  Q  vdd pp ww='5'
Xn3  Q   Qn gnd nn ww='5'
Xp4  Q   Qn vdd pp ww='5'
Xn5  bff wl Qn  nn ww='5'
Xn6  btt wl Q   nn ww='5'
.ends mem1



.subckt decode2 o11 o10 o01 o00 di1 di0 df1 df0
Xn11 o11 di1 di0 nnd2 size=10
Xn10 o10 di1 df0 nnd2 size=10
Xn01 o01 df1 di0 nnd2 size=10
Xn00 o00 df1 df0 nnd2 size=10
.ends


.subckt decode_nor16 k1111 k1110 k1101 k1100 k1011 k1010 k1001 k1000 k0111 k0101

.ends

.subckt decode_nnd16

.ends


.subckt decode_16and1

.ends decode_16and1


.subckt dmux256 o255 o223 0012 o001 dt7 dt6 dt5 d4 dt3 dt1 dt0

.ends dmux256






