

* File includes subcircuits and technology definitions
.include ./SRAM_bits.cir


*this cell emulates load from SRAM cells,
* Number refers to the load from than number of cells
.subckt memLoad ttt fff number=254
Xnt ttt gnd dead nn ww='number*5'
Xnf fff gnd dead nn ww='number*5'
.ends memLoad




*********begin: topLevel*****

* Parameters
.global gnd vdd
.param gnd=0


*********begin: topLevel*****
.param per = 5ns
.param lw=500
.param wirew=3


*DC supplies
vdd vdd 0 'supply'
Xclok clk               dat1 period='0.5*per' total=1 duty=0.5 sz=120
Xrdwr rdw               dat1 period='per' start='per' total=2 duty=1
*Vrdw rdw 0 'supply'
Xbit  ad0               dat1 period='per' start='per' total=3 duty=1
*Vdii dii 0 '0'
Xacc acc                dat1 period='per' start='per+10ps' total=2 duty=1

*
Xwr bt0 bf0 dii rdw clk write1
Xw0 bt0 bt1 bf0 bf1     wire_dual len='lw' wid='wirew'
Xla bt1 bf1 ope         mem1 m=1
Xmd bt1 bf1             memLoad number =254

Xw1 bt1 bt2 bf1 bf2     wire_dual len='lw' wid='wirew'
Xrd bt2 bf2 dot rdw clk read1

Xde ope ad0 clk decModel size=100



.tran 1p 25n






