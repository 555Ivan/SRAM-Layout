

* File includes subcircuits and technology definitions
.include ./SRAM_bits.cir



.subckt SRAM a7 a6 a5 a4 a3 a2 a1 a0
+            w7 w6 w5 w4 w3 w2 w1 w0
+            r7 r6 r5 r4 r3 r2 r1 r0
+            rw ck

*SRAM cell
Xw w7 w6 w5 w4 w3 w2 w1 w0
+   it7 it6 it5 it4 it3 it2 it1 it0
+   if7 if6 if5 if4 if3 if2 if1 if0
+   rw clk write

* this is a single 8-bit word cell
* need 256
Xm it7 it6 it5 it4 it3 it2 it1 it0
+   if7 if6 if5 if4 if3 if2 if1 if0
+   ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0
+   of7 of6 of5 of4 of3 of2 of1 of0
+   acc mem8


Xr r7 r6 r5 r4 r3 r2 r1 r0
+   ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0
+   of7 of6 of5 of4 of3 of2 of1 of0
+   rw clk read

* demux only outputs eight choices for simplicity
Xd c7 c6 c5 c4 c3 c2 c1 c0
+	a7 a6 a5 a4 a3 a2 a1 a0 demux256
.ends SRAM


* address is a[7:0]
* only 8 of 256 combinations exported here,
.subckt demux256 c7 c6 c5 c4 c3 c2 c1 c0
+	             a7 a6 a5 a4 a3 a2 a1 a0
.ends demux256


.subckt write di7 di6 di5 di4 di3 di2 di1 di0
+              bt7 bt6 bt5 bt4 bt3 bt2 bt1 bt0
+              bf7 bf6 bf5 bf4 bf3 bf2 bf1 bf0
+              rw clk
* connect 8 read circuits here
X0 bt0 bf0 di0 rw clk write1
.ends write


.subckt mem8  it7 it6 it5 it4 it3 it2 it1 it0
+              if7 if6 if5 if4 if3 if2 if1 if0
+              ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0
+              of7 of6 of5 of4 of3 of2 of1 of0
+              acc wid='wid' len='len'
X7 it7 if7 ot7 of7 ac mem1 wid='wid' len='len'
X6 it6 if6 ot6 of6 ac mem1 wid='wid' len='len'
X5 it5 if5 ot5 of5 ac mem1 wid='wid' len='len'
X4 it4 if4 ot4 of4 ac mem1 wid='wid' len='len'
X3 it3 if3 ot3 of3 ac mem1 wid='wid' len='len'
X2 it2 if2 ot2 of2 ac mem1 wid='wid' len='len'
X1 it1 if1 ot1 of1 ac mem1 wid='wid' len='len'
X0 it0 if0 ot0 of0 ac mem1 wid='wid' len='len'
.ends mem8

.subckt mem1 it if ot of ac wid=10 len=10
Xwrt it ot wire wid='wid' len='len'
Xwrf if of wire wid='wid' len='len'
xpst it ac tt  nn ww=5
xpsf if ac ff  nn ww=5
Xpif tt ff vdd pp ww=5
xpit ff tt vdd pp ww=5
Xnit tt ff gnd nn ww=5
xnif ff tt gnd nn ww=5
.ends mem1


.subckt read ot7 ot6 ot5 ot4 ot3 ot2 ot1 ot0
+             bt7 bt6 bt5 bt4 bt3 bt2 bt1 bt0
+             bf7 bf6 bf5 bf4 bf3 bf2 bf1 bf0
+            rw clk
* connect 8 read circuits here
X1 ot0 bt0 bf0 rw clk read1
.ends read



* Parameters
.global gnd vdd
.param gnd=0


*********begin: topLevel*****
.param per = 1ns


*DC supplies
vdd vdd 0 'supply'
Xclok clk               dat1 per='0.5*per' total=1 dut=0.5 sz=120
Xrdwr rdw               dat1 per='per' start='per' total=6 duty=1


* This register (reg8)  passes the address bits generated by (dat8)
Xgad8 gd7 gd6 gd5 gd4 gd3 gd2 gd1 gd0     dat8 per='per' start='per'
Xadd8 ad7 ad6 ad5 ad4 ad3 ad2 ad1 ad0
+     gd7 gd6 gd5 gd4 gd3 gd2 gd1 gd0 clk reg8

* This register (reg8)  passes the bits for
*writing into the SRAM that are generated by (dat8)
Xgwr8 di7 di6 di5 di4 di3 di2 di1 di0     dat8 per='per' start='per'
Xrdw8 wr7 wr6 wr5 wr4 wr3 wr2 wr1 wr0
+     di7 di6 di5 di4 di3 di2 di1 di0 clk reg8

*This register consumes data from the SRAM
Xred8 oo7 oo6 oo5 oo4 oo3 oo2 oo1 oo0
+    do7 do6 do5 do4 do3 do2 do1 do0 clk  reg8

*This is an 256 element x 8bit word SRAM
Xsram ad7 ad6 ad5 ad4 ad3 ad2 ad1 ad0
+      wr7 wr6 wr5 wr4 wr3 wr2 wr1 wr0
+      o7 do6 do5 do4 do3 do2 do1 do0
+      rdw clk sram



.tran 1p 28n
*Below is the format for stepping a parameter while re-running a simulation
*.step param ddd 1.93ns 2.07n 0.007n


* measurement statement

*.meas ivdd find i(vdd) at=1.8n
*.meas thresh find v(thr) at=1.8n
*.meas del1 trig v(n1) val='0.5*supply' rise =2 targ v(n1) val='0.5*supply'   rise=3
*.meas de param = 'del10/70'
*.meas rtime  trig v(n2) val= '0.1 * supply' rise = 2 targ v(n2) val = '0.9*supply' rise =2
*.meas ftime  trig v(n2) val= '0.9 * supply' fall = 2 targ v(n2) val = '0.1*supply' fall =2





